module Example4( output logic    out
               , input  logic    a
               , input  logic[2] bc
               );

   nand n1(out, a, ab[1]);

endmodule;
