primitive collect
  ( output logic o
  , input  logic a
  , input  logic b
  );

   assign o = a;
   assign o = b;

endprimitive; // collect
