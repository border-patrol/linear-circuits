module Example1( input  logic a
               , input  logic b
               , output logic c);

   wire logic as (o,i);

   and(c,a,b);

endmodule;
