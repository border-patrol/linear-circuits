module Example6( output logic    o
               , input  logic    i
               );

   assign o = i;

endmodule;
