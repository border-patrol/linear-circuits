module BVEdgesGood ( output logic      o
                  , input  logic[1:0] i);

   and a(o,i[1],i[0]);

endmodule; // BVEdges
