module Mux ( output logic a
           , input  logic b
           , input  logic c
           , input  logic d);

   mux m(a,b,c,d);

endmodule; // BVEdges
