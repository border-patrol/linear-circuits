primitive split
  ( output logic a
  , output logic b
  , input logic i
  );

   assign a = i;
   assign b = i;

endprimitive; // split
