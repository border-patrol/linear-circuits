module SimpleAssignment( output logic    o
              , input  logic    i
              );

   assign o = i;

endmodule;
