module Example6( input  logic    a
               , input  logic    b
               , output logic[2] c
               );

   merge(c, a, b);

endmodule;
